module divider4
